-- Vhdl test bench created from schematic D:\digitalLogic_slides\random\prj1\test4.sch - Mon Jan 29 22:04:59 2018
--
-- Notes: 
-- 1) This testbench template has been automatically generated using types
-- std_logic and std_logic_vector for the ports of the unit under test.
-- Xilinx recommends that these types always be used for the top-level
-- I/O of a design in order to guarantee that the testbench will bind
-- correctly to the timing (post-route) simulation model.
-- 2) To use this template as your testbench, change the filename to any
-- name of your choice with the extension .vhd, and use the "Source->Add"
-- menu in Project Navigator to import the testbench. Then
-- edit the user defined section below, adding code to generate the 
-- stimulus for your design.
--
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
LIBRARY UNISIM;
USE UNISIM.Vcomponents.ALL;
ENTITY test4_test4_sch_tb IS
END test4_test4_sch_tb;
ARCHITECTURE behavioral OF test4_test4_sch_tb IS 

   COMPONENT test4
   PORT( clear	:	IN	STD_LOGIC; 
          clk	:	IN	STD_LOGIC; 
          c	:	OUT	STD_LOGIC_VECTOR (7 DOWNTO 0); 
          roll	:	IN	STD_LOGIC; 
			 user	:	OUT	STD_LOGIC;
			 m :	OUT	STD_LOGIC;
			 Win0 :	OUT	STD_LOGIC;
			 Win1 :	OUT	STD_LOGIC;
			 stop	:	IN	STD_LOGIC; 
          B	:	OUT	STD_LOGIC_VECTOR (3 DOWNTO 0); 
          S	:	OUT	STD_LOGIC_VECTOR (7 DOWNTO 0);
			 Score0	:	OUT	STD_LOGIC_VECTOR (7 DOWNTO 0);
			  Score1	:	OUT	STD_LOGIC_VECTOR (7 DOWNTO 0));
   END COMPONENT;

   SIGNAL clear	:	STD_LOGIC;
   SIGNAL clk	:	STD_LOGIC;
	SIGNAL stop	:	STD_LOGIC;
	SIGNAL user	:	STD_LOGIC;
   SIGNAL c	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
   SIGNAL roll	:	STD_LOGIC;
	SIGNAL m	:	STD_LOGIC;
	SIGNAL Win0	:	STD_LOGIC;
	SIGNAL Win1	:	STD_LOGIC;
   SIGNAL B	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
   SIGNAL S	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL Score0	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL Score1	:	STD_LOGIC_VECTOR (7 DOWNTO 0);	

BEGIN

   UUT: test4 PORT MAP(
		clear => clear, 
		clk => clk, 
		c => c, 
		roll => roll, 
		B => B, 
		S => S,
		user => user,
		Score0 => Score0,
		Score1 => Score1,
		stop => stop,
		m => m,
		Win0 =>Win0,
		Win1 =>Win1
	);

-- *** Test Bench - User Defined Section ***
   tb : PROCESS
   BEGIN
	
	clk <='1';
	clear <='1';
	roll <='0';
	stop <='0';
	wait for 25 ns;
	clk<='0';
	clear<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll <='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop <='1'; 
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<= '1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	stop<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	stop<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	stop<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	stop<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	stop<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	stop<='0';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='1';
	wait for 25 ns;
	clk<='1';
	wait for 25 ns;
	clk<='0';
	roll<='0';
	wait for 25 ns;
	clk<='1';
	roll<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	roll<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	stop<='1';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;
	clk<='1';
	stop<='0';
	wait for 25 ns;
	clk<='0';
	wait for 25 ns;	
      WAIT; -- will wait forever
   END PROCESS;
-- *** End Test Bench - User Defined Section ***

END;
